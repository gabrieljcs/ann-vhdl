../../ann-vhdl/src/network_test.vhd
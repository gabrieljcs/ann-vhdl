../src/network.vhd
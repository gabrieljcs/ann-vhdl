../src/neuron.vhd
../src/act_func.vhd
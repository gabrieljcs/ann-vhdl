../src/types.vhd
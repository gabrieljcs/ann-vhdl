../src/network_test_tb.vhd